module mod7_fsm (
    input   clk,
    input   rst_n,
    input   data_in,

    output reg [2:0]    data_out
);
    
endmodule