module clk_div (
    input  rst_n,
    input  clk_100mhz,
    output clk_100hz,
    output clk_25mhz
);



endmodule
